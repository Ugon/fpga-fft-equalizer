library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fft_twiddle_factors_16 is
	type arr is array (0 to 7) of signed(23 downto 0);
	
	constant tw_size: integer := 24;

	constant re_16: arr := (
		0 => "011111111111111111111111", --one
		1 => "011101100100000110101111",
		2 => "010110101000001001111010",
		3 => "001100001111101111000101",
		4 => "000000000000000000000000",
		5 => "110011110000010000111011",
		6 => "101001010111110110000110",
		7 => "100010011011111001010001");

	constant im_16: arr := (
		0 => "000000000000000000000000",
		1 => "001100001111101111000101",
		2 => "010110101000001001111010",
		3 => "011101100100000110101111",
		4 => "011111111111111111111111", --one
		5 => "011101100100000110101111",
		6 => "010110101000001001111010",
		7 => "001100001111101111000101");

end;