library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fft_twiddle_factors_256 is
	constant tw_size:           integer := 24;
	constant tw_array_size_exp: integer := 8;
	
	type arr is array (0 to 127) of signed(tw_size - 1 downto 0);

	constant re_256: arr := (
		0 =>"011111111111111111111111",  --one 24-bit approximation
		1 =>"011111111111011000100010",
		2 =>"011111111101100010001000",
		3 =>"011111111010011100110111",
		4 =>"011111110110001000110111",
		5 =>"011111110000100110010010",
		6 =>"011111101001110101010110",
		7 =>"011111100001110110010100",
		8 =>"011111011000101001011111",
		9 =>"011111001110001111001111",
		10 =>"011111000010100111111100",
		11 =>"011110110101110100000100",
		12 =>"011110100111110100000101",
		13 =>"011110011000101000100100",
		14 =>"011110001000010010000100",
		15 =>"011101110110110001001111",
		16 =>"011101100100000110101111",
		17 =>"011101010000010011010011",
		18 =>"011100111011010111101100",
		19 =>"011100100101010100101101",
		20 =>"011100001110001011001100",
		21 =>"011011110101111100000011",
		22 =>"011011011100101000001101",
		23 =>"011011000010010000101001",
		24 =>"011010100110110110011001",
		25 =>"011010001010011010011111",
		26 =>"011001101100111110000001",
		27 =>"011001001110100010001001",
		28 =>"011000101111001000000010",
		29 =>"011000001110110000111000",
		30 =>"010111101101011101111101",
		31 =>"010111001011010000100001",
		32 =>"010110101000001001111010",
		33 =>"010110000100001011011101",
		34 =>"010101011111010110100101",
		35 =>"010100111001101100101011",
		36 =>"010100010011001111001101",
		37 =>"010011101011111111101001",
		38 =>"010011000011111111100000",
		39 =>"010010011011010000010101",
		40 =>"010001110001110011101101",
		41 =>"010001000111101011001101",
		42 =>"010000011100111000011110",
		43 =>"001111110001011101001010",
		44 =>"001111000101011010111010",
		45 =>"001110011000110011011101",
		46 =>"001101101011101000100000",
		47 =>"001100111101111011110011",
		48 =>"001100001111101111000101",
		49 =>"001011100001000100001010",
		50 =>"001010110001111100110101",
		51 =>"001010000010011010111001",
		52 =>"001001010010100000001100",
		53 =>"001000100010001110100101",
		54 =>"000111110001100111111001",
		55 =>"000111000000101110000010",
		56 =>"000110001111100010111000",
		57 =>"000101011110001000010100",
		58 =>"000100101100100000010000",
		59 =>"000011111010101100100111",
		60 =>"000011001000101111010011",
		61 =>"000010010110101010010000",
		62 =>"000001100100011111011001",
		63 =>"000000110010010000101011",
		64 =>"000000000000000000000000",
		65 =>"111111001101101111010101",
		66 =>"111110011011100000100111",
		67 =>"111101101001010101110000",
		68 =>"111100110111010000101101",
		69 =>"111100000101010011011001",
		70 =>"111011010011011111110000",
		71 =>"111010100001110111101100",
		72 =>"111001110000011101001000",
		73 =>"111000111111010001111110",
		74 =>"111000001110011000000111",
		75 =>"110111011101110001011011",
		76 =>"110110101101011111110100",
		77 =>"110101111101100101000111",
		78 =>"110101001110000011001011",
		79 =>"110100011110111011110110",
		80 =>"110011110000010000111011",
		81 =>"110011000010000100001101",
		82 =>"110010010100010111100000",
		83 =>"110001100111001100100011",
		84 =>"110000111010100101000110",
		85 =>"110000001110100010110110",
		86 =>"101111100011000111100010",
		87 =>"101110111000010100110011",
		88 =>"101110001110001100010011",
		89 =>"101101100100101111101011",
		90 =>"101100111100000000100000",
		91 =>"101100010100000000010111",
		92 =>"101011101100110000110011",
		93 =>"101011000110010011010101",
		94 =>"101010100000101001011011",
		95 =>"101001111011110100100011",
		96 =>"101001010111110110000110",
		97 =>"101000110100101111011111",
		98 =>"101000010010100010000011",
		99 =>"100111110001001111001000",
		100 =>"100111010000110111111110",
		101 =>"100110110001011101110111",
		102 =>"100110010011000001111111",
		103 =>"100101110101100101100001",
		104 =>"100101011001001001100111",
		105 =>"100100111101101111010111",
		106 =>"100100100011010111110011",
		107 =>"100100001010000011111101",
		108 =>"100011110001110100110100",
		109 =>"100011011010101011010011",
		110 =>"100011000100101000010100",
		111 =>"100010101111101100101101",
		112 =>"100010011011111001010001",
		113 =>"100010001001001110110001",
		114 =>"100001110111101101111100",
		115 =>"100001100111010111011100",
		116 =>"100001011000001011111011",
		117 =>"100001001010001011111100",
		118 =>"100000111101011000000100",
		119 =>"100000110001110000110001",
		120 =>"100000100111010110100001",
		121 =>"100000011110001001101100",
		122 =>"100000010110001010101010",
		123 =>"100000001111011001101110",
		124 =>"100000001001110111001001",
		125 =>"100000000101100011001001",
		126 =>"100000000010011101111000",
		127 =>"100000000000100111011110");

	constant im_256: arr := (
		0 =>"000000000000000000000000",
		1 =>"000000110010010000101011",
		2 =>"000001100100011111011001",
		3 =>"000010010110101010010000",
		4 =>"000011001000101111010011",
		5 =>"000011111010101100100111",
		6 =>"000100101100100000010000",
		7 =>"000101011110001000010100",
		8 =>"000110001111100010111000",
		9 =>"000111000000101110000010",
		10 =>"000111110001100111111001",
		11 =>"001000100010001110100101",
		12 =>"001001010010100000001100",
		13 =>"001010000010011010111001",
		14 =>"001010110001111100110101",
		15 =>"001011100001000100001010",
		16 =>"001100001111101111000101",
		17 =>"001100111101111011110011",
		18 =>"001101101011101000100000",
		19 =>"001110011000110011011101",
		20 =>"001111000101011010111010",
		21 =>"001111110001011101001010",
		22 =>"010000011100111000011110",
		23 =>"010001000111101011001101",
		24 =>"010001110001110011101101",
		25 =>"010010011011010000010101",
		26 =>"010011000011111111100000",
		27 =>"010011101011111111101001",
		28 =>"010100010011001111001101",
		29 =>"010100111001101100101011",
		30 =>"010101011111010110100101",
		31 =>"010110000100001011011101",
		32 =>"010110101000001001111010",
		33 =>"010111001011010000100001",
		34 =>"010111101101011101111101",
		35 =>"011000001110110000111000",
		36 =>"011000101111001000000010",
		37 =>"011001001110100010001001",
		38 =>"011001101100111110000001",
		39 =>"011010001010011010011111",
		40 =>"011010100110110110011001",
		41 =>"011011000010010000101001",
		42 =>"011011011100101000001101",
		43 =>"011011110101111100000011",
		44 =>"011100001110001011001100",
		45 =>"011100100101010100101101",
		46 =>"011100111011010111101100",
		47 =>"011101010000010011010011",
		48 =>"011101100100000110101111",
		49 =>"011101110110110001001111",
		50 =>"011110001000010010000100",
		51 =>"011110011000101000100100",
		52 =>"011110100111110100000101",
		53 =>"011110110101110100000100",
		54 =>"011111000010100111111100",
		55 =>"011111001110001111001111",
		56 =>"011111011000101001011111",
		57 =>"011111100001110110010100",
		58 =>"011111101001110101010110",
		59 =>"011111110000100110010010",
		60 =>"011111110110001000110111",
		61 =>"011111111010011100110111",
		62 =>"011111111101100010001000",
		63 =>"011111111111011000100010",
		64 =>"011111111111111111111111",  --one 24-bit approximation
		65 =>"011111111111011000100010",
		66 =>"011111111101100010001000",
		67 =>"011111111010011100110111",
		68 =>"011111110110001000110111",
		69 =>"011111110000100110010010",
		70 =>"011111101001110101010110",
		71 =>"011111100001110110010100",
		72 =>"011111011000101001011111",
		73 =>"011111001110001111001111",
		74 =>"011111000010100111111100",
		75 =>"011110110101110100000100",
		76 =>"011110100111110100000101",
		77 =>"011110011000101000100100",
		78 =>"011110001000010010000100",
		79 =>"011101110110110001001111",
		80 =>"011101100100000110101111",
		81 =>"011101010000010011010011",
		82 =>"011100111011010111101100",
		83 =>"011100100101010100101101",
		84 =>"011100001110001011001100",
		85 =>"011011110101111100000011",
		86 =>"011011011100101000001101",
		87 =>"011011000010010000101001",
		88 =>"011010100110110110011001",
		89 =>"011010001010011010011111",
		90 =>"011001101100111110000001",
		91 =>"011001001110100010001001",
		92 =>"011000101111001000000010",
		93 =>"011000001110110000111000",
		94 =>"010111101101011101111101",
		95 =>"010111001011010000100001",
		96 =>"010110101000001001111010",
		97 =>"010110000100001011011101",
		98 =>"010101011111010110100101",
		99 =>"010100111001101100101011",
		100 =>"010100010011001111001101",
		101 =>"010011101011111111101001",
		102 =>"010011000011111111100000",
		103 =>"010010011011010000010101",
		104 =>"010001110001110011101101",
		105 =>"010001000111101011001101",
		106 =>"010000011100111000011110",
		107 =>"001111110001011101001010",
		108 =>"001111000101011010111010",
		109 =>"001110011000110011011101",
		110 =>"001101101011101000100000",
		111 =>"001100111101111011110011",
		112 =>"001100001111101111000101",
		113 =>"001011100001000100001010",
		114 =>"001010110001111100110101",
		115 =>"001010000010011010111001",
		116 =>"001001010010100000001100",
		117 =>"001000100010001110100101",
		118 =>"000111110001100111111001",
		119 =>"000111000000101110000010",
		120 =>"000110001111100010111000",
		121 =>"000101011110001000010100",
		122 =>"000100101100100000010000",
		123 =>"000011111010101100100111",
		124 =>"000011001000101111010011",
		125 =>"000010010110101010010000",
		126 =>"000001100100011111011001",
		127 =>"000000110010010000101011");

end;