library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fft_twiddle_factors_64 is
	constant tw_size:           integer := 16;
	constant tw_array_size_exp: integer := 6;
	
	type arr is array (0 to 2**(tw_array_size_exp - 1) - 1) of signed(tw_size - 1 downto 0);

	constant re_64: arr := (
		0 =>  "0111111111111111", --'one' 16-bit approximation
		1 =>  "0111111101100010",
		2 =>  "0111110110001010",
		3 =>  "0111101001111101",
		4 =>  "0111011001000010",
		5 =>  "0111000011100011",
		6 =>  "0110101001101110",
		7 =>  "0110001011110010",
		8 =>  "0101101010000010",
		9 =>  "0101000100110100",
		10 => "0100011100011101",
		11 => "0011110001010111",
		12 => "0011000011111100",
		13 => "0010010100101000",
		14 => "0001100011111001",
		15 => "0000110010001100",
		16 => "0000000000000000",
		17 => "1111001101110100",
		18 => "1110011100000111",
		19 => "1101101011011000",
		20 => "1100111100000100",
		21 => "1100001110101001",
		22 => "1011100011100011",
		23 => "1010111011001100",
		24 => "1010010101111110",
		25 => "1001110100001110",
		26 => "1001010110010010",
		27 => "1000111100011101",
		28 => "1000100110111110",
		29 => "1000010110000011",
		30 => "1000001001110110",
		31 => "1000000010011110");

	constant im_64: arr := (
		0 =>  "0000000000000000",
		1 =>  "0000110010001100",
		2 =>  "0001100011111001",
		3 =>  "0010010100101000",
		4 =>  "0011000011111100",
		5 =>  "0011110001010111",
		6 =>  "0100011100011101",
		7 =>  "0101000100110100",
		8 =>  "0101101010000010",
		9 =>  "0110001011110010",
		10 => "0110101001101110",
		11 => "0111000011100011",
		12 => "0111011001000010",
		13 => "0111101001111101",
		14 => "0111110110001010",
		15 => "0111111101100010",
		16 => "0111111111111111", --'one' 16-bit approximation
		17 => "0111111101100010",
		18 => "0111110110001010",
		19 => "0111101001111101",
		20 => "0111011001000010",
		21 => "0111000011100011",
		22 => "0110101001101110",
		23 => "0110001011110010",
		24 => "0101101010000010",
		25 => "0101000100110100",
		26 => "0100011100011101",
		27 => "0011110001010111",
		28 => "0011000011111100",
		29 => "0010010100101000",
		30 => "0001100011111001",
		31 => "0000110010001100");

end;